module bcd7seg(b,h);
  input [3:0] b;
  output reg [7:0] h;
  
  always @(b) begin
    case (b)
        4'b0000 : h = 8'b01000000;
        4'b0001 : h = 8'b01111001;
        4'b0010 : h = 8'b00100100;
        4'b0011 : h = 8'b00110000;
        4'b0100 : h = 8'b00011001;
        4'b0101 : h = 8'b00010010;
        4'b0110 : h = 8'b00000010;
        4'b0111 : h = 8'b01111000;
        4'b1000 : h = 8'b00000000;
        4'b1001 : h = 8'b00010000;
        4'b1010 : h = 8'b00001000;
        4'b1011 : h = 8'b00000011;
        4'b1100 : h = 8'b01000110;
        4'b1101 : h = 8'b00100001;
        4'b1110 : h = 8'b00000110;
        4'b1111 : h = 8'b00001110;
    endcase
  end
endmodule
